module IDU();
endmodule;
