module IFU #(
)(
);

endmodule;
