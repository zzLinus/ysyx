module EXU();
endmodule;
