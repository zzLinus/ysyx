	// verilator_coverage annotation
	module top(
 000021		input clk,
%000002	  input rst
	);
	
	endmodule;
	
