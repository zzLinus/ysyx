module lookup_table(
	input [7:0] key_code,
	output [7:0] ascii_code
);

endmodule
