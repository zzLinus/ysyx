module IFU();
endmodule;
