module adder (

)
