// module shift_register(
// 	input clk,
// 	input data,
// 	output out_q
// );
//
// endmodule
